module _and(input A, B, output C);

assign C= A&B;


endmodule 