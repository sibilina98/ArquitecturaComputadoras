//1.Definicion del modulo y sus entradas y salidas
module _and(input A, input B, output C );
//2. Declarar señales/elementos internos
//NA
//3.Comportamiento del modulo
//  (asifnaciones, instanicas, conexiones)
assign C = A&B; 

endmodule
//https://github.com/sibilina98/ArquitecturaComputadoras.git 